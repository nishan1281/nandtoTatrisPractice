<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-5.31661,-1.67645,68.9834,-89.8765</PageViewport>
<gate>
<ID>2</ID>
<type>AA_TOGGLE</type>
<position>6.5,-28</position>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>18.5,-28</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>30,-28</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_TOGGLE</type>
<position>40,-28</position>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>20</ID>
<type>AA_AND4</type>
<position>60,-34</position>
<input>
<ID>IN_0</ID>14 </input>
<input>
<ID>IN_1</ID>9 </input>
<input>
<ID>IN_2</ID>8 </input>
<input>
<ID>IN_3</ID>13 </input>
<output>
<ID>OUT</ID>1 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_AND4</type>
<position>60,-45</position>
<input>
<ID>IN_0</ID>14 </input>
<input>
<ID>IN_1</ID>10 </input>
<input>
<ID>IN_2</ID>8 </input>
<input>
<ID>IN_3</ID>13 </input>
<output>
<ID>OUT</ID>2 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>24</ID>
<type>AA_AND4</type>
<position>60,-56</position>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>11 </input>
<input>
<ID>IN_2</ID>8 </input>
<input>
<ID>IN_3</ID>13 </input>
<output>
<ID>OUT</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>26</ID>
<type>AA_AND4</type>
<position>60.5,-66.5</position>
<input>
<ID>IN_0</ID>11 </input>
<input>
<ID>IN_1</ID>10 </input>
<input>
<ID>IN_2</ID>8 </input>
<input>
<ID>IN_3</ID>13 </input>
<output>
<ID>OUT</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>30</ID>
<type>AE_SMALL_INVERTER</type>
<position>12.5,-28</position>
<input>
<ID>IN_0</ID>11 </input>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>32</ID>
<type>AE_SMALL_INVERTER</type>
<position>24,-28</position>
<input>
<ID>IN_0</ID>10 </input>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>34</ID>
<type>GA_LED</type>
<position>64,-34</position>
<input>
<ID>N_in0</ID>1 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>36</ID>
<type>GA_LED</type>
<position>64,-45</position>
<input>
<ID>N_in0</ID>2 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>38</ID>
<type>GA_LED</type>
<position>64,-56</position>
<input>
<ID>N_in0</ID>3 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>40</ID>
<type>GA_LED</type>
<position>65,-66.5</position>
<input>
<ID>N_in0</ID>4 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63,-34,63,-34</points>
<connection>
<GID>34</GID>
<name>N_in0</name></connection>
<connection>
<GID>20</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63,-45,63,-45</points>
<connection>
<GID>36</GID>
<name>N_in0</name></connection>
<connection>
<GID>22</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63,-56,63,-56</points>
<connection>
<GID>38</GID>
<name>N_in0</name></connection>
<connection>
<GID>24</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>63.5,-66.5,64,-66.5</points>
<connection>
<GID>40</GID>
<name>N_in0</name></connection>
<connection>
<GID>26</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,-67.5,36,-28</points>
<intersection>-67.5 2</intersection>
<intersection>-57 4</intersection>
<intersection>-46 6</intersection>
<intersection>-35 8</intersection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32,-28,36,-28</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>36 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>36,-67.5,57.5,-67.5</points>
<connection>
<GID>26</GID>
<name>IN_2</name></connection>
<intersection>36 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>36,-57,57,-57</points>
<connection>
<GID>24</GID>
<name>IN_2</name></connection>
<intersection>36 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>36,-46,57,-46</points>
<connection>
<GID>22</GID>
<name>IN_2</name></connection>
<intersection>36 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>36,-35,57,-35</points>
<connection>
<GID>20</GID>
<name>IN_2</name></connection>
<intersection>36 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26,-33,57,-33</points>
<connection>
<GID>20</GID>
<name>IN_1</name></connection>
<intersection>26 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>26,-53,26,-28</points>
<connection>
<GID>32</GID>
<name>OUT_0</name></connection>
<intersection>-53 5</intersection>
<intersection>-33 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>26,-53,57,-53</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>26 3</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>21,-44,57,-44</points>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<intersection>21 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>21,-65.5,21,-28</points>
<intersection>-65.5 7</intersection>
<intersection>-44 1</intersection>
<intersection>-28 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>20.5,-28,22,-28</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<connection>
<GID>32</GID>
<name>IN_0</name></connection>
<intersection>21 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>21,-65.5,57.5,-65.5</points>
<connection>
<GID>26</GID>
<name>IN_1</name></connection>
<intersection>21 3</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>8.5,-28,10.5,-28</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>9.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>9.5,-63.5,9.5,-28</points>
<intersection>-63.5 7</intersection>
<intersection>-55 5</intersection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>9.5,-55,57,-55</points>
<connection>
<GID>24</GID>
<name>IN_1</name></connection>
<intersection>9.5 4</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>9.5,-63.5,57.5,-63.5</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>9.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47,-69.5,47,-28</points>
<intersection>-69.5 2</intersection>
<intersection>-59 5</intersection>
<intersection>-48 4</intersection>
<intersection>-37 3</intersection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>42,-28,47,-28</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>47 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>47,-69.5,57.5,-69.5</points>
<connection>
<GID>26</GID>
<name>IN_3</name></connection>
<intersection>47 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>47,-37,57,-37</points>
<connection>
<GID>20</GID>
<name>IN_3</name></connection>
<intersection>47 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>47,-48,57,-48</points>
<connection>
<GID>22</GID>
<name>IN_3</name></connection>
<intersection>47 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>47,-59,57,-59</points>
<connection>
<GID>24</GID>
<name>IN_3</name></connection>
<intersection>47 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>14.5,-31,57,-31</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>14.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>14.5,-42,14.5,-28</points>
<connection>
<GID>30</GID>
<name>OUT_0</name></connection>
<intersection>-42 5</intersection>
<intersection>-31 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>14.5,-42,57,-42</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>14.5 3</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,74.3,-88.2</PageViewport></page 1>
<page 2>
<PageViewport>0,0,74.3,-88.2</PageViewport></page 2>
<page 3>
<PageViewport>0,0,74.3,-88.2</PageViewport></page 3>
<page 4>
<PageViewport>0,0,74.3,-88.2</PageViewport></page 4>
<page 5>
<PageViewport>0,0,74.3,-88.2</PageViewport></page 5>
<page 6>
<PageViewport>0,0,74.3,-88.2</PageViewport></page 6>
<page 7>
<PageViewport>0,0,74.3,-88.2</PageViewport></page 7>
<page 8>
<PageViewport>0,0,74.3,-88.2</PageViewport></page 8>
<page 9>
<PageViewport>0,0,74.3,-88.2</PageViewport></page 9></circuit>